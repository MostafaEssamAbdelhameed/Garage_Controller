`timescale 1ns / 1ps


module door_tb();
parameter clk_period= 20;
reg clk_tb=0;
always #(clk_period/2) clk_tb = ~clk_tb;

///////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////
reg UP_max_tb , activate_tb , DN_max_tb , rst_tb;
wire UP_m_tb , DN_m_tb;

door DUT (  .UP_max(UP_max_tb),
            .activate(activate_tb),
            .DN_max(DN_max_tb),
            .rst(rst_tb),
            .clk(clk_tb),
            .UP_m(UP_m_tb),
            .DN_m(DN_m_tb)
            );
///////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////            
initial begin 
   // do_op(UP_max,Activate,DN_max);

    initialize();
    do_op(1,1,0);
    do_op(0,1,1);
    do_op(1,0,0);
    
    #(2*clk_period)

    $stop;

end            
///////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////
task initialize ;
    begin
        rst_tb=0;
        activate_tb = 0;
    end
endtask
///////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////
task reset;
    begin
    rst_tb = 1;
    #(clk_period)
    rst_tb=0;
    #(clk_period)
    rst_tb = 1;
    end
endtask
///////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////
task do_op;
    input up_max , activate , dn_max ;
    begin 
        reset();
       // #(clk_period)
        activate_tb = activate;
        UP_max_tb=up_max;
        DN_max_tb = dn_max;
        #(clk_period)

        $display("Sensor up = %d ",UP_max_tb,
                 "Sensor Down = %d ",DN_max_tb,
                 "so set Up motor = %d and Down Motor = %d",UP_m_tb,DN_m_tb);
        UP_max_tb=0;
        DN_max_tb=0;                 
    end
endtask
///////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////
endmodule
